// Time-stamp: <2021-05-07 16:34:15 kmodi>

program top;

  initial begin
    $hello;
    $bye;

    $finish;
  end

endprogram : top
