// Time-stamp: <2021-05-07 12:27:51 kmodi>

program top;

  initial begin
    $hello;
    $finish;
  end

endprogram : top
