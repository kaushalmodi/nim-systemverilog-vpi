// Time-stamp: <2021-05-19 09:13:03 kmodi>

program top;

  initial begin
    $bye;

    $finish;
  end

endprogram : top
