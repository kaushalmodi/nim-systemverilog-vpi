orig/tb.sv