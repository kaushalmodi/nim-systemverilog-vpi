orig/vlab_probes_pkg.sv